module ISM(
	input logic CLK,
	input logic RESET,
	input logic transition1.
	input logic transition2,
	input logic calculating,
	output logic [1:0] state
);



endmodule
