'define img_width 640
'define img_height 480
module fractal_calc(


);
begin

	real real_var, cpx_var;
	string color_var;



	get_color rgbgen();

	always_comb
	begin
		for ()
		begin
			for ()
			begin
				
			end
		end
	end
	
endmodule
