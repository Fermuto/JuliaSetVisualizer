module ISM(

);
begin

endmodule
