// jsv_sdram.v

// Generated using ACDS version 19.1 670

`timescale 1 ps / 1 ps
module jsv_sdram (
		input  wire [22:0] bridge_0_ext_address,     // bridge_0_ext.address
		input  wire [1:0]  bridge_0_ext_byte_enable, //             .byte_enable
		input  wire        bridge_0_ext_read,        //             .read
		input  wire        bridge_0_ext_write,       //             .write
		input  wire [15:0] bridge_0_ext_write_data,  //             .write_data
		output wire        bridge_0_ext_acknowledge, //             .acknowledge
		output wire [15:0] bridge_0_ext_read_data,   //             .read_data
		input  wire        clk_clk,                  //          clk.clk
		input  wire        reset_reset_n,            //        reset.reset_n
		output wire        sdram_clk_clk,            //    sdram_clk.clk
		output wire [11:0] sdram_wire_addr,          //   sdram_wire.addr
		output wire        sdram_wire_ba,            //             .ba
		output wire        sdram_wire_cas_n,         //             .cas_n
		output wire        sdram_wire_cke,           //             .cke
		output wire        sdram_wire_cs_n,          //             .cs_n
		inout  wire [15:0] sdram_wire_dq,            //             .dq
		output wire [1:0]  sdram_wire_dqm,           //             .dqm
		output wire        sdram_wire_ras_n,         //             .ras_n
		output wire        sdram_wire_we_n           //             .we_n
	);

	wire         sdram_pll_c0_clk;                                // sdram_pll:c0 -> [bitmap_sdram:clk, mm_interconnect_0:sdram_pll_c0_clk, rst_controller:clk]
	wire  [15:0] bridge_0_avalon_master_readdata;                 // mm_interconnect_0:bridge_0_avalon_master_readdata -> bridge_0:avalon_readdata
	wire         bridge_0_avalon_master_waitrequest;              // mm_interconnect_0:bridge_0_avalon_master_waitrequest -> bridge_0:avalon_waitrequest
	wire   [1:0] bridge_0_avalon_master_byteenable;               // bridge_0:avalon_byteenable -> mm_interconnect_0:bridge_0_avalon_master_byteenable
	wire         bridge_0_avalon_master_read;                     // bridge_0:avalon_read -> mm_interconnect_0:bridge_0_avalon_master_read
	wire  [22:0] bridge_0_avalon_master_address;                  // bridge_0:avalon_address -> mm_interconnect_0:bridge_0_avalon_master_address
	wire         bridge_0_avalon_master_write;                    // bridge_0:avalon_write -> mm_interconnect_0:bridge_0_avalon_master_write
	wire  [15:0] bridge_0_avalon_master_writedata;                // bridge_0:avalon_writedata -> mm_interconnect_0:bridge_0_avalon_master_writedata
	wire  [31:0] mm_interconnect_0_sdram_pll_pll_slave_readdata;  // sdram_pll:readdata -> mm_interconnect_0:sdram_pll_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_sdram_pll_pll_slave_address;   // mm_interconnect_0:sdram_pll_pll_slave_address -> sdram_pll:address
	wire         mm_interconnect_0_sdram_pll_pll_slave_read;      // mm_interconnect_0:sdram_pll_pll_slave_read -> sdram_pll:read
	wire         mm_interconnect_0_sdram_pll_pll_slave_write;     // mm_interconnect_0:sdram_pll_pll_slave_write -> sdram_pll:write
	wire  [31:0] mm_interconnect_0_sdram_pll_pll_slave_writedata; // mm_interconnect_0:sdram_pll_pll_slave_writedata -> sdram_pll:writedata
	wire         mm_interconnect_0_bitmap_sdram_s1_chipselect;    // mm_interconnect_0:bitmap_sdram_s1_chipselect -> bitmap_sdram:az_cs
	wire  [15:0] mm_interconnect_0_bitmap_sdram_s1_readdata;      // bitmap_sdram:za_data -> mm_interconnect_0:bitmap_sdram_s1_readdata
	wire         mm_interconnect_0_bitmap_sdram_s1_waitrequest;   // bitmap_sdram:za_waitrequest -> mm_interconnect_0:bitmap_sdram_s1_waitrequest
	wire  [20:0] mm_interconnect_0_bitmap_sdram_s1_address;       // mm_interconnect_0:bitmap_sdram_s1_address -> bitmap_sdram:az_addr
	wire         mm_interconnect_0_bitmap_sdram_s1_read;          // mm_interconnect_0:bitmap_sdram_s1_read -> bitmap_sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_bitmap_sdram_s1_byteenable;    // mm_interconnect_0:bitmap_sdram_s1_byteenable -> bitmap_sdram:az_be_n
	wire         mm_interconnect_0_bitmap_sdram_s1_readdatavalid; // bitmap_sdram:za_valid -> mm_interconnect_0:bitmap_sdram_s1_readdatavalid
	wire         mm_interconnect_0_bitmap_sdram_s1_write;         // mm_interconnect_0:bitmap_sdram_s1_write -> bitmap_sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_bitmap_sdram_s1_writedata;     // mm_interconnect_0:bitmap_sdram_s1_writedata -> bitmap_sdram:az_data
	wire         rst_controller_reset_out_reset;                  // rst_controller:reset_out -> [bitmap_sdram:reset_n, mm_interconnect_0:bitmap_sdram_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset;              // rst_controller_001:reset_out -> [bridge_0:reset, mm_interconnect_0:bridge_0_reset_reset_bridge_in_reset_reset, sdram_pll:reset]

	jsv_sdram_bitmap_sdram bitmap_sdram (
		.clk            (sdram_pll_c0_clk),                                //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                 // reset.reset_n
		.az_addr        (mm_interconnect_0_bitmap_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_bitmap_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_bitmap_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_bitmap_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_bitmap_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_bitmap_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_bitmap_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_bitmap_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_bitmap_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                                 //  wire.export
		.zs_ba          (sdram_wire_ba),                                   //      .export
		.zs_cas_n       (sdram_wire_cas_n),                                //      .export
		.zs_cke         (sdram_wire_cke),                                  //      .export
		.zs_cs_n        (sdram_wire_cs_n),                                 //      .export
		.zs_dq          (sdram_wire_dq),                                   //      .export
		.zs_dqm         (sdram_wire_dqm),                                  //      .export
		.zs_ras_n       (sdram_wire_ras_n),                                //      .export
		.zs_we_n        (sdram_wire_we_n)                                  //      .export
	);

	jsv_sdram_bridge_0 bridge_0 (
		.clk                (clk_clk),                            //                clk.clk
		.reset              (rst_controller_001_reset_out_reset), //              reset.reset
		.avalon_readdata    (bridge_0_avalon_master_readdata),    //      avalon_master.readdata
		.avalon_waitrequest (bridge_0_avalon_master_waitrequest), //                   .waitrequest
		.avalon_byteenable  (bridge_0_avalon_master_byteenable),  //                   .byteenable
		.avalon_read        (bridge_0_avalon_master_read),        //                   .read
		.avalon_write       (bridge_0_avalon_master_write),       //                   .write
		.avalon_writedata   (bridge_0_avalon_master_writedata),   //                   .writedata
		.avalon_address     (bridge_0_avalon_master_address),     //                   .address
		.address            (bridge_0_ext_address),               // external_interface.export
		.byte_enable        (bridge_0_ext_byte_enable),           //                   .export
		.read               (bridge_0_ext_read),                  //                   .export
		.write              (bridge_0_ext_write),                 //                   .export
		.write_data         (bridge_0_ext_write_data),            //                   .export
		.acknowledge        (bridge_0_ext_acknowledge),           //                   .export
		.read_data          (bridge_0_ext_read_data)              //                   .export
	);

	jsv_sdram_sdram_pll sdram_pll (
		.clk                (clk_clk),                                         //       inclk_interface.clk
		.reset              (rst_controller_001_reset_out_reset),              // inclk_interface_reset.reset
		.read               (mm_interconnect_0_sdram_pll_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_sdram_pll_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_sdram_pll_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_sdram_pll_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_sdram_pll_pll_slave_writedata), //                      .writedata
		.c0                 (sdram_pll_c0_clk),                                //                    c0.clk
		.c1                 (sdram_clk_clk),                                   //                    c1.clk
		.scandone           (),                                                //           (terminated)
		.scandataout        (),                                                //           (terminated)
		.c2                 (),                                                //           (terminated)
		.c3                 (),                                                //           (terminated)
		.c4                 (),                                                //           (terminated)
		.areset             (1'b0),                                            //           (terminated)
		.locked             (),                                                //           (terminated)
		.phasedone          (),                                                //           (terminated)
		.phasecounterselect (3'b000),                                          //           (terminated)
		.phaseupdown        (1'b0),                                            //           (terminated)
		.phasestep          (1'b0),                                            //           (terminated)
		.scanclk            (1'b0),                                            //           (terminated)
		.scanclkena         (1'b0),                                            //           (terminated)
		.scandata           (1'b0),                                            //           (terminated)
		.configupdate       (1'b0)                                             //           (terminated)
	);

	jsv_sdram_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                  (clk_clk),                                         //                                clk_0_clk.clk
		.sdram_pll_c0_clk                               (sdram_pll_c0_clk),                                //                             sdram_pll_c0.clk
		.bitmap_sdram_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                  // bitmap_sdram_reset_reset_bridge_in_reset.reset
		.bridge_0_reset_reset_bridge_in_reset_reset     (rst_controller_001_reset_out_reset),              //     bridge_0_reset_reset_bridge_in_reset.reset
		.bridge_0_avalon_master_address                 (bridge_0_avalon_master_address),                  //                   bridge_0_avalon_master.address
		.bridge_0_avalon_master_waitrequest             (bridge_0_avalon_master_waitrequest),              //                                         .waitrequest
		.bridge_0_avalon_master_byteenable              (bridge_0_avalon_master_byteenable),               //                                         .byteenable
		.bridge_0_avalon_master_read                    (bridge_0_avalon_master_read),                     //                                         .read
		.bridge_0_avalon_master_readdata                (bridge_0_avalon_master_readdata),                 //                                         .readdata
		.bridge_0_avalon_master_write                   (bridge_0_avalon_master_write),                    //                                         .write
		.bridge_0_avalon_master_writedata               (bridge_0_avalon_master_writedata),                //                                         .writedata
		.bitmap_sdram_s1_address                        (mm_interconnect_0_bitmap_sdram_s1_address),       //                          bitmap_sdram_s1.address
		.bitmap_sdram_s1_write                          (mm_interconnect_0_bitmap_sdram_s1_write),         //                                         .write
		.bitmap_sdram_s1_read                           (mm_interconnect_0_bitmap_sdram_s1_read),          //                                         .read
		.bitmap_sdram_s1_readdata                       (mm_interconnect_0_bitmap_sdram_s1_readdata),      //                                         .readdata
		.bitmap_sdram_s1_writedata                      (mm_interconnect_0_bitmap_sdram_s1_writedata),     //                                         .writedata
		.bitmap_sdram_s1_byteenable                     (mm_interconnect_0_bitmap_sdram_s1_byteenable),    //                                         .byteenable
		.bitmap_sdram_s1_readdatavalid                  (mm_interconnect_0_bitmap_sdram_s1_readdatavalid), //                                         .readdatavalid
		.bitmap_sdram_s1_waitrequest                    (mm_interconnect_0_bitmap_sdram_s1_waitrequest),   //                                         .waitrequest
		.bitmap_sdram_s1_chipselect                     (mm_interconnect_0_bitmap_sdram_s1_chipselect),    //                                         .chipselect
		.sdram_pll_pll_slave_address                    (mm_interconnect_0_sdram_pll_pll_slave_address),   //                      sdram_pll_pll_slave.address
		.sdram_pll_pll_slave_write                      (mm_interconnect_0_sdram_pll_pll_slave_write),     //                                         .write
		.sdram_pll_pll_slave_read                       (mm_interconnect_0_sdram_pll_pll_slave_read),      //                                         .read
		.sdram_pll_pll_slave_readdata                   (mm_interconnect_0_sdram_pll_pll_slave_readdata),  //                                         .readdata
		.sdram_pll_pll_slave_writedata                  (mm_interconnect_0_sdram_pll_pll_slave_writedata)  //                                         .writedata
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (sdram_pll_c0_clk),               //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
