module visualizer_top(

);
begin



endmodule
