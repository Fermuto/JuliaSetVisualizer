module naturallog(
    input int x,
    output logic [31:0] y
);
    always_comb
    begin
        case (x)
            1: y = 32'b0000000000000000_0000000000000000;
            2: y = 32'b0000000000000000_1011000101110010;
            3: y = 32'b0000000000000001_0001100100111110;
            4: y = 32'b0000000000000001_0110001011100100;
            5: y = 32'b0000000000000001_1001110000000100;
            6: y = 32'b0000000000000001_1100101010110000;
            7: y = 32'b0000000000000001_1111001000100111;
            8: y = 32'b0000000000000010_0001010001010110;
            9: y = 32'b0000000000000010_0011001001111101;
            10: y = 32'b0000000000000010_0100110101110110;
            11: y = 32'b0000000000000010_0110010111011100;
            12: y = 32'b0000000000000010_0111110000100010;
            13: y = 32'b0000000000000010_1001000010100000;
            14: y = 32'b0000000000000010_1010001110011001;
            15: y = 32'b0000000000000010_1011010101000010;
            16: y = 32'b0000000000000010_1100010111001000;
            17: y = 32'b0000000000000010_1101010101001101;
            18: y = 32'b0000000000000010_1110001111101111;
            19: y = 32'b0000000000000010_1111000111000110;
            20: y = 32'b0000000000000010_1111111011101000;
            21: y = 32'b0000000000000011_0000101101100101;
            22: y = 32'b0000000000000011_0001011101001110;
            23: y = 32'b0000000000000011_0010001010101111;
            24: y = 32'b0000000000000011_0010110110010100;
            25: y = 32'b0000000000000011_0011100000001000;
            26: y = 32'b0000000000000011_0100001000010010;
            27: y = 32'b0000000000000011_0100101110111011;
            28: y = 32'b0000000000000011_0101010100001011;
            29: y = 32'b0000000000000011_0101111000000111;
            30: y = 32'b0000000000000011_0110011010110100;
            31: y = 32'b0000000000000011_0110111100011001;
            32: y = 32'b0000000000000011_0111011100111010;
            33: y = 32'b0000000000000011_0111111100011011;
            34: y = 32'b0000000000000011_1000011010111111;
            35: y = 32'b0000000000000011_1000111000101011;
            36: y = 32'b0000000000000011_1001010101100001;
            37: y = 32'b0000000000000011_1001110001100101;
            38: y = 32'b0000000000000011_1010001100111000;
            39: y = 32'b0000000000000011_1010100111011111;
            40: y = 32'b0000000000000011_1011000001011010;
            41: y = 32'b0000000000000011_1011011010101100;
            42: y = 32'b0000000000000011_1011110011010111;
            43: y = 32'b0000000000000011_1100001011011110;
            44: y = 32'b0000000000000011_1100100011000000;
            45: y = 32'b0000000000000011_1100111010000001;
            46: y = 32'b0000000000000011_1101010000100001;
            47: y = 32'b0000000000000011_1101100110100011;
            48: y = 32'b0000000000000011_1101111100000111;
            49: y = 32'b0000000000000011_1110010001001110;
            50: y = 32'b0000000000000011_1110100101111010;
            51: y = 32'b0000000000000011_1110111010001100;
            52: y = 32'b0000000000000011_1111001110000100;
            53: y = 32'b0000000000000011_1111100001100101;
            54: y = 32'b0000000000000011_1111110100101110;
            55: y = 32'b0000000000000100_0000000111100000;
            56: y = 32'b0000000000000100_0000011001111101;
            57: y = 32'b0000000000000100_0000101100000101;
            58: y = 32'b0000000000000100_0000111101111001;
            59: y = 32'b0000000000000100_0001001111011001;
            60: y = 32'b0000000000000100_0001100000100110;
            61: y = 32'b0000000000000100_0001110001100010;
            62: y = 32'b0000000000000100_0010000010001011;
            63: y = 32'b0000000000000100_0010010010100100;
            64: y = 32'b0000000000000100_0010100010101100;
            65: y = 32'b0000000000000100_0010110010100100;
            66: y = 32'b0000000000000100_0011000010001101;
            67: y = 32'b0000000000000100_0011010001100110;
            68: y = 32'b0000000000000100_0011100000110001;
            69: y = 32'b0000000000000100_0011101111101110;
            70: y = 32'b0000000000000100_0011111110011101;
            71: y = 32'b0000000000000100_0100001100111110;
            72: y = 32'b0000000000000100_0100011011010011;
            73: y = 32'b0000000000000100_0100101001011011;
            74: y = 32'b0000000000000100_0100110111010111;
            75: y = 32'b0000000000000100_0101000101000110;
            76: y = 32'b0000000000000100_0101010010101010;
            77: y = 32'b0000000000000100_0101100000000011;
            78: y = 32'b0000000000000100_0101101101010001;
            79: y = 32'b0000000000000100_0101111010010100;
            80: y = 32'b0000000000000100_0110000111001100;
            81: y = 32'b0000000000000100_0110010011111010;
            82: y = 32'b0000000000000100_0110100000011110;
            83: y = 32'b0000000000000100_0110101100111001;
            84: y = 32'b0000000000000100_0110111001001010;
            85: y = 32'b0000000000000100_0111000101010001;
            86: y = 32'b0000000000000100_0111010001010000;
            87: y = 32'b0000000000000100_0111011101000101;
            88: y = 32'b0000000000000100_0111101000110010;
            89: y = 32'b0000000000000100_0111110100010111;
            90: y = 32'b0000000000000100_0111111111110011;
            91: y = 32'b0000000000000100_1000001011000111;
            92: y = 32'b0000000000000100_1000010110010011;
            93: y = 32'b0000000000000100_1000100001011000;
            94: y = 32'b0000000000000100_1000101100010101;
            95: y = 32'b0000000000000100_1000110111001010;
            96: y = 32'b0000000000000100_1001000001111001;
            97: y = 32'b0000000000000100_1001001100100000;
            98: y = 32'b0000000000000100_1001010111000000;
            99: y = 32'b0000000000000100_1001100001011001;
            100: y = 32'b0000000000000100_1001101011101100;
            101: y = 32'b0000000000000100_1001110101111000;
				default: y = 32'b0000000000000000_0000000000000000;
        endcase
    end
endmodule