module fractal_calc(


);
begin

real real_var, cpx_var;
string color_var;

endmodule
